library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_ARITH.all;
use IEEE.STD_LOGIC_UNSIGNED.all;

-- Created from etherhm2.bin
-- On 9/14/2023

entity etherhm2 is
	port (
	addr: in std_logic_vector(11 downto 0);
	clk: in std_logic;
	din: in std_logic_vector(23 downto 0);
	dout: out std_logic_vector(23 downto 0);
	we: in std_logic);
end etherhm2;

architecture syn of etherhm2 is
   type ram_type is array (0 to 4095) of std_logic_vector(23 downto 0);
   signal RAM : ram_type := 
   (
   x"000000", x"000000", x"000000", x"010000", x"8F0000",
   x"10025A", x"10039C", x"1003FF", x"100318", x"100239",
   x"40013A", x"330000", x"40012C", x"330011", x"010000",
   x"B00079", x"200013", x"010001", x"B00079", x"4B0000",
   x"B0007A", x"4000B0", x"330019", x"400031", x"33000C",
   x"40007C", x"B00150", x"01017F", x"850000", x"1000A0",
   x"32000C", x"010180", x"850000", x"000000", x"000000",
   x"010800", x"060000", x"E90006", x"320040", x"010806",
   x"060000", x"E90006", x"32002E", x"000000", x"000000",
   x"20000C", x"4000A8", x"E90013", x"33000C", x"4000A9",
   x"E90014", x"33000C", x"0104B6", x"840000", x"010806",
   x"060000", x"B000B6", x"010040", x"B000B4", x"100419",
   x"10018C", x"10019B", x"10010F", x"20000C", x"4000A8",
   x"E9000F", x"330046", x"4000A9", x"E90010", x"32004E",
   x"4000A8", x"5000AC", x"E9000F", x"33000C", x"4000A9",
   x"5000AD", x"E90010", x"33000C", x"49000B", x"E0008F",
   x"70008D", x"320059", x"49000B", x"E00090", x"70008D",
   x"32006E", x"000000", x"000000", x"20000C", x"010180",
   x"840000", x"4000B1", x"B000B4", x"010800", x"060000",
   x"B000B6", x"10018C", x"1001D7", x"1001F2", x"01FFF2",
   x"C080B1", x"014001", x"060000", x"B8000B", x"000000",
   x"4000B1", x"060000", x"B80008", x"10010F", x"20000C",
   x"490012", x"E000D8", x"33000C", x"490013", x"060000",
   x"E00088", x"0B0000", x"B000DC", x"0104CB", x"840000",
   x"010195", x"850000", x"40007C", x"B00151", x"2004A9",
   x"B000B4", x"32000A", x"010001", x"C08134", x"0104B6",
   x"840000", x"010180", x"850000", x"010008", x"C080B4",
   x"010800", x"060000", x"B000B6", x"10018C", x"1001D7",
   x"1001F9", x"4000B4", x"060000", x"B80013", x"010014",
   x"C080B4", x"014011", x"060000", x"B8000B", x"4000B4",
   x"060000", x"B80008", x"01000E", x"C080B4", x"40007C",
   x"B00152", x"10010F", x"40007C", x"B00153", x"20000A",
   x"B0003C", x"4000B0", x"3300B8", x"000000", x"01C092",
   x"100156", x"40009F", x"B0009E", x"01C092", x"100143",
   x"012000", x"70009F", x"3200FA", x"010000", x"B0009E",
   x"013090", x"100143", x"01309C", x"100156", x"01FF00",
   x"70009F", x"060000", x"B000B0", x"320104", x"000000",
   x"01FFFF", x"C080B0", x"01307C", x"100156", x"018000",
   x"70009F", x"320100", x"010017", x"70009F", x"330100",
   x"013C00", x"70009F", x"330100", x"000000", x"01C07E",
   x"100156", x"010FFF", x"70009F", x"B000B1", x"B000B2",
   x"320100", x"014000", x"B0009E", x"01C086", x"100143",
   x"010238", x"B0009E", x"01C082", x"100143", x"10016C",
   x"10016C", x"10016C", x"C00083", x"70008E", x"B000B2",
   x"E000B9", x"3C0100", x"B00041", x"400045", x"000000",
   x"000000", x"000000", x"000000", x"400041", x"B90000",
   x"400045", x"000000", x"000000", x"000000", x"000000",
   x"400041", x"B90001", x"01FFFC", x"C080B2", x"890002",
   x"3300DF", x"000000", x"010230", x"B0009E", x"01C082",
   x"100143", x"012800", x"B0009E", x"013090", x"100143",
   x"010001", x"C08130", x"01FFFA", x"C080B1", x"B0003D",
   x"280000", x"010231", x"B0009E", x"01C082", x"100143",
   x"012800", x"B0009E", x"013090", x"100143", x"010008",
   x"50812C", x"010001", x"C08132", x"010000", x"B0003D",
   x"280000", x"B0003E", x"4000B4", x"C00083", x"70008E",
   x"B000B5", x"E000B8", x"3C013D", x"010238", x"B0009E",
   x"01C082", x"100143", x"018000", x"100174", x"4000B4",
   x"100174", x"B00051", x"480000", x"B00030", x"B00059",
   x"000000", x"000000", x"000000", x"480001", x"B00051",
   x"B00030", x"B00059", x"000000", x"880002", x"000000",
   x"000000", x"B00051", x"01FFFC", x"C080B5", x"33011F",
   x"010230", x"B0009E", x"01C082", x"100143", x"010001",
   x"B0009E", x"013080", x"100143", x"010001", x"C08133",
   x"B0003F", x"280000", x"010001", x"C08135", x"010010",
   x"50812C", x"B0003F", x"280000", x"B00030", x"B00053",
   x"B0005B", x"000000", x"000000", x"000000", x"000000",
   x"B00053", x"40009E", x"B00030", x"B00051", x"B00059",
   x"000000", x"000000", x"000000", x"000000", x"B00051",
   x"B00040", x"280000", x"B00030", x"B00053", x"B0005B",
   x"000000", x"000000", x"000000", x"000000", x"B00053",
   x"B00041", x"B00045", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"400030",
   x"B0009F", x"000000", x"B00041", x"280000", x"400041",
   x"400045", x"000000", x"000000", x"000000", x"000000",
   x"400041", x"280000", x"B00030", x"B00051", x"B00059",
   x"000000", x"000000", x"000000", x"000000", x"B00051",
   x"280000", x"4000A5", x"B80000", x"4000A6", x"B80001",
   x"4000A7", x"B80002", x"4000A2", x"B80003", x"4000A3",
   x"B80004", x"4000A4", x"B80005", x"4000B6", x"B80006",
   x"280000", x"490003", x"B80000", x"490004", x"B80001",
   x"490005", x"B80002", x"4000A2", x"B80003", x"4000A3",
   x"B80004", x"4000A4", x"B80005", x"4000B6", x"B80006",
   x"280000", x"010001", x"060000", x"B80007", x"010800",
   x"060000", x"B80008", x"010604", x"060000", x"B80009",
   x"010002", x"060000", x"B8000A", x"4000A2", x"B8000B",
   x"4000A3", x"B8000C", x"4000A4", x"B8000D", x"4000A8",
   x"B8000E", x"4000A9", x"B8000F", x"49000B", x"B80010",
   x"49000C", x"B80011", x"49000D", x"B80012", x"49000E",
   x"B80013", x"49000F", x"B80014", x"280000", x"014500",
   x"060000", x"B80007", x"010000", x"060000", x"B80008",
   x"010000", x"060000", x"B80009", x"014000", x"060000",
   x"B8000A", x"014011", x"060000", x"B8000B", x"010000",
   x"060000", x"B8000C", x"4000A8", x"B8000D", x"4000AA",
   x"B8000E", x"4000AE", x"B8000F", x"4000AF", x"B80010",
   x"280000", x"014500", x"060000", x"B80007", x"010000",
   x"060000", x"B80008", x"010000", x"060000", x"B80009",
   x"014000", x"060000", x"B8000A", x"014011", x"060000",
   x"B8000B", x"010000", x"060000", x"B8000C", x"49000D",
   x"B8000F", x"49000E", x"B80010", x"4000A8", x"B8000D",
   x"4000A9", x"B8000E", x"280000", x"010000", x"060000",
   x"B80011", x"010000", x"060000", x"B80012", x"280000",
   x"490011", x"B80012", x"4000D8", x"B80011", x"010000",
   x"060000", x"B80014", x"280000", x"010044", x"060000",
   x"B80011", x"010043", x"060000", x"B80012", x"010134",
   x"060000", x"B80013", x"010000", x"060000", x"B80014",
   x"280000", x"010101", x"060000", x"B80015", x"010600",
   x"060000", x"B80016", x"4000BC", x"B80017", x"4000BD",
   x"B80018", x"010001", x"060000", x"B80019", x"018000",
   x"060000", x"B8001A", x"4000A8", x"B8001B", x"4000A9",
   x"B8001C", x"010000", x"060000", x"B8001D", x"010000",
   x"060000", x"B8001E", x"4000AE", x"B8001F", x"4000AF",
   x"B80020", x"010000", x"060000", x"B80021", x"010000",
   x"060000", x"B80022", x"4000A2", x"B80023", x"4000A3",
   x"B80024", x"4000A4", x"B80025", x"280000", x"01FFFF",
   x"B0007B", x"011111", x"B0007A", x"010064", x"100450",
   x"012222", x"B0007A", x"010064", x"100450", x"014444",
   x"B0007A", x"010064", x"100450", x"018888", x"B0007A",
   x"010064", x"100450", x"014444", x"B0007A", x"010064",
   x"100450", x"012222", x"B0007A", x"010064", x"100450",
   x"011111", x"B0007A", x"010064", x"100450", x"400136",
   x"B0007B", x"280000", x"100429", x"015A00", x"B00154",
   x"015A01", x"B0015C", x"015A02", x"B0011C", x"015A03",
   x"B00100", x"015A04", x"B00165", x"015A06", x"B00124",
   x"015A07", x"B0013C", x"016F48", x"B00158", x"017473",
   x"B00159", x"016F4D", x"B0015A", x"013274", x"B0015B",
   x"01534B", x"B00160", x"01385A", x"B00161", x"013538",
   x"B00162", x"010031", x"B00163", x"017445", x"B00120",
   x"016568", x"B00121", x"014572", x"B00122", x"015045",
   x"B00123", x"015046", x"B00104", x"014147", x"B00105",
   x"016C46", x"B00106", x"016873", x"B00107", x"016954",
   x"B00169", x"01656D", x"B0016A", x"017372", x"B0016B",
   x"010000", x"B0016C", x"01424C", x"B00128", x"013150",
   x"B00129", x"015236", x"B0012A", x"010057", x"B0012B",
   x"01424C", x"B00140", x"013150", x"B00141", x"015236",
   x"B00142", x"01004F", x"B00143", x"010130", x"870000",
   x"010008", x"B00137", x"010003", x"B0014C", x"010012",
   x"B0014D", x"010001", x"B00081", x"010002", x"B00082",
   x"010003", x"B00083", x"010004", x"B00084", x"010005",
   x"B00085", x"010006", x"B00086", x"010007", x"B00087",
   x"010008", x"B00088", x"010010", x"B0008A", x"01000F",
   x"B00091", x"018104", x"B00155", x"010010", x"B00156",
   x"018102", x"B0015D", x"010008", x"B0015E", x"018E02",
   x"B0011D", x"010007", x"B0011E", x"018F04", x"B00101",
   x"018200", x"B00102", x"018202", x"B00166", x"010004",
   x"B00167", x"018202", x"B00125", x"010004", x"B00126",
   x"010202", x"B0013D", x"010004", x"B0013E", x"0100FF",
   x"B0008C", x"01FF00", x"B0008D", x"01FFFC", x"B0008E",
   x"010100", x"B0008F", x"011100", x"B00090", x"010400",
   x"B00092", x"010800", x"B00093", x"010C00", x"B00094",
   x"011000", x"B00095", x"011800", x"B00097", x"011C00",
   x"B00098", x"010100", x"B00099", x"010200", x"B0009A",
   x"01000F", x"B000EA", x"010060", x"060000", x"B000A2",
   x"011B10", x"060000", x"B000A3", x"010000", x"060000",
   x"B000A4", x"01FF00", x"060000", x"B000A5", x"010000",
   x"060000", x"B000A6", x"010000", x"060000", x"B000A7",
   x"016A2D", x"060000", x"B000D8", x"010044", x"060000",
   x"B000DA", x"010600", x"B000B9", x"010600", x"B000B8",
   x"0104B1", x"B000BB", x"0107FB", x"B000BA", x"01FFFF",
   x"B0007D", x"280000", x"01FFFF", x"060000", x"B000AA",
   x"01FF00", x"060000", x"B000AB", x"010003", x"70003F",
   x"B0014E", x"E00081", x"320328", x"E00081", x"320341",
   x"000000", x"000000", x"20038F", x"010011", x"B000D5",
   x"100812", x"4000D4", x"060000", x"B000A8", x"010010",
   x"B000D5", x"100812", x"4000D4", x"060000", x"B000A9",
   x"010013", x"B000D5", x"100812", x"4000D4", x"060000",
   x"B000AA", x"010012", x"B000D5", x"100812", x"4000D4",
   x"060000", x"B000AB", x"200395", x"10043B", x"4000D0",
   x"B000BC", x"4000D1", x"B000BD", x"0104B6", x"840000",
   x"010148", x"B000B4", x"100419", x"010800", x"060000",
   x"B000B6", x"01FFFF", x"B000AE", x"B000AF", x"B000A5",
   x"B000A6", x"B000A7", x"010000", x"B000A8", x"B000A9",
   x"014011", x"060000", x"B8000B", x"10017D", x"1001BC",
   x"4000B4", x"060000", x"B80008", x"01000E", x"C080B4",
   x"100201", x"10020E", x"10010F", x"0103E8", x"B0009D",
   x"010001", x"100450", x"01FFFF", x"C0809D", x"320341",
   x"4000B0", x"33036F", x"400031", x"330366", x"000000",
   x"000000", x"01017F", x"850000", x"1000A0", x"320366",
   x"010180", x"850000", x"000000", x"000000", x"010800",
   x"060000", x"E90006", x"330366", x"49000B", x"E00090",
   x"70008D", x"330366", x"490012", x"E000DA", x"330366",
   x"490017", x"E000BC", x"330366", x"490018", x"E000BD",
   x"330366", x"49001D", x"B000A8", x"49001E", x"B000A9",
   x"200395", x"01C0A8", x"060000", x"B000A8", x"010179",
   x"060000", x"B000A9", x"01FFFF", x"6000AA", x"B000AC",
   x"01FFFF", x"6000AB", x"B000AD", x"280000", x"000000",
   x"010000", x"B00032", x"01000A", x"100450", x"010001",
   x"B00032", x"01000A", x"100450", x"010001", x"B0009E",
   x"01C026", x"100143", x"01000A", x"100450", x"010000",
   x"B0009E", x"01C026", x"100143", x"01000A", x"100450",
   x"013014", x"100156", x"40009F", x"70008C", x"B0009E",
   x"013014", x"100143", x"40009E", x"060000", x"B000A2",
   x"01C012", x"100156", x"40009F", x"060000", x"B000A3",
   x"013010", x"100156", x"40009F", x"060000", x"B000A4",
   x"014000", x"B0009E", x"013084", x"100143", x"0101EE",
   x"B0009E", x"013070", x"100143", x"014000", x"B0009E",
   x"01C086", x"100143", x"010001", x"B0009E", x"01309C",
   x"100143", x"017CE0", x"B0009E", x"013074", x"100143",
   x"010016", x"B0009E", x"01C076", x"100143", x"010230",
   x"B0009E", x"01C082", x"100143", x"0120FF", x"B0009E",
   x"01C0F6", x"100143", x"01FFFF", x"B0009E", x"01C092",
   x"100143", x"012800", x"B0009E", x"013090", x"100143",
   x"0101EF", x"B0009E", x"013070", x"100143", x"017CE1",
   x"B0009E", x"013074", x"100143", x"4000A4", x"B000CC",
   x"B000CD", x"4000A3", x"B000CE", x"B000CF", x"000000",
   x"000000", x"000000", x"280000", x"010008", x"B000D5",
   x"010000", x"860000", x"100812", x"4000D4", x"BA0144",
   x"010001", x"C080D5", x"820000", x"E00087", x"3C040E",
   x"8A0001", x"000000", x"200403", x"010014", x"B000D5",
   x"100812", x"4000D4", x"B00136", x"B0007B", x"1008E3",
   x"010004", x"C000E6", x"508102", x"280000", x"0B0000",
   x"B0009C", x"0104B6", x"860000", x"010000", x"BA0000",
   x"000000", x"000000", x"000000", x"01FFFF", x"8A0001",
   x"C0809C", x"33041D", x"000000", x"000000", x"280000",
   x"010080", x"860000", x"010000", x"BA0000", x"000000",
   x"000000", x"000000", x"8A0001", x"820000", x"040000",
   x"040000", x"040000", x"040000", x"040000", x"3C042B",
   x"000000", x"000000", x"280000", x"019069", x"A000CC",
   x"C000CD", x"B000CC", x"080000", x"D00080", x"B000CD",
   x"014650", x"A000CE", x"C000CF", x"B000CE", x"080000",
   x"D00080", x"B000CF", x"4000CE", x"B000D0", x"000000",
   x"4000CF", x"C000CD", x"B000D1", x"280000", x"B000BE",
   x"0137CE", x"B000BF", x"000000", x"000000", x"01FFFF",
   x"C080BF", x"000000", x"000000", x"330455", x"01FFFF",
   x"C080BE", x"330451", x"000000", x"000000", x"280000",
   x"011100", x"B00068", x"01FFFF", x"B00060", x"B00061",
   x"B0006D", x"000000", x"000000", x"000000", x"011104",
   x"B00068", x"01FFFF", x"B00060", x"B00061", x"B0006D",
   x"000000", x"000000", x"000000", x"011108", x"B00068",
   x"01FFFF", x"B00060", x"B00061", x"B0006D", x"000000",
   x"000000", x"000000", x"01110C", x"B00068", x"01FFFF",
   x"B00060", x"B00061", x"B0006D", x"000000", x"000000",
   x"000000", x"011000", x"B00068", x"010000", x"B00060",
   x"B00061", x"B0006D", x"000000", x"000000", x"000000",
   x"011004", x"B00068", x"010000", x"B00060", x"B00061",
   x"B0006D", x"000000", x"000000", x"000000", x"011008",
   x"B00068", x"010000", x"B00060", x"B00061", x"B0006D",
   x"000000", x"000000", x"000000", x"01100C", x"B00068",
   x"010000", x"B00060", x"B00061", x"B0006D", x"000000",
   x"000000", x"000000", x"280000", x"810000", x"C000DC",
   x"B000DD", x"800000", x"B000DE", x"490000", x"B000DF",
   x"000000", x"890001", x"01007F", x"7000DF", x"3204F6",
   x"B0009B", x"013C00", x"7000DF", x"330511", x"010300",
   x"7000DF", x"E0009A", x"3304F6", x"014000", x"7000DF",
   x"3204C4", x"490000", x"B00157", x"890001", x"2004C5",
   x"400157", x"B00068", x"018000", x"7000DF", x"3304DA",
   x"B0006C", x"800000", x"E000BA", x"3C04FE", x"4000DF",
   x"B0006E", x"400060", x"B80000", x"400061", x"B80001",
   x"01FFFF", x"C0809B", x"880002", x"3304C9", x"400068",
   x"B00157", x"2004EB", x"490000", x"B00060", x"490001",
   x"B00061", x"810000", x"E000BB", x"3C04FE", x"B0006D",
   x"890002", x"4000DF", x"B0006E", x"01FFFF", x"C0809B",
   x"3304DA", x"000000", x"400068", x"B00157", x"810000",
   x"E000DD", x"3804AE", x"010001", x"C08131", x"010000",
   x"B00139", x"800000", x"E000DE", x"040000", x"20007D",
   x"010001", x"50812C", x"01FFFF", x"E0012D", x"32050D",
   x"010001", x"C0812D", x"20050D", x"010002", x"50812C",
   x"01FFFF", x"E0012E", x"32050D", x"010001", x"C0812E",
   x"20050D", x"010004", x"50812C", x"01FFFF", x"E0012F",
   x"32050D", x"010001", x"C0812F", x"010000", x"B00139",
   x"8F0000", x"20007D", x"011C00", x"7000DF", x"E00095",
   x"3205E1", x"011C00", x"7000DF", x"E00092", x"3206AA",
   x"011C00", x"7000DF", x"E00093", x"320707", x"011C00",
   x"7000DF", x"E00094", x"320768", x"011C00", x"7000DF",
   x"E00098", x"32052F", x"011C00", x"7000DF", x"E00097",
   x"320569", x"011C00", x"7000DF", x"320697", x"000000",
   x"000000", x"2004F6", x"012000", x"7000DF", x"330556",
   x"010300", x"7000DF", x"E00099", x"3304F6", x"014000",
   x"7000DF", x"32053D", x"490000", x"B0013F", x"890001",
   x"20053F", x"000000", x"40013F", x"0B0000", x"860000",
   x"018000", x"7000DF", x"330506", x"820000", x"E0008A",
   x"3C04FE", x"4A0144", x"B80000", x"010080", x"7000DF",
   x"32054F", x"010002", x"C0813F", x"8A0001", x"01FFFF",
   x"C0809B", x"880001", x"330544", x"000000", x"000000",
   x"2004EB", x"1007E1", x"820000", x"E00088", x"3C04FE",
   x"4A013C", x"B80000", x"010080", x"7000DF", x"320562",
   x"010002", x"C080E2", x"8A0001", x"01FFFF", x"C0809B",
   x"880001", x"330557", x"000000", x"000000", x"2004EB",
   x"012000", x"7000DF", x"3305CE", x"010300", x"7000DF",
   x"E00099", x"3304F6", x"014000", x"7000DF", x"320577",
   x"490000", x"B00127", x"890001", x"200578", x"400127",
   x"0B0000", x"860000", x"018000", x"7000DF", x"3305A5",
   x"820000", x"E0008A", x"3C04FE", x"820000", x"E000EA",
   x"330596", x"010001", x"B00022", x"000000", x"000000",
   x"010001", x"B00021", x"000000", x"000000", x"000000",
   x"010000", x"B00021", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"400020", x"B80000", x"200598",
   x"4A012C", x"B80000", x"010080", x"7000DF", x"32059E",
   x"010002", x"C08127", x"8A0001", x"01FFFF", x"C0809B",
   x"880001", x"33057D", x"000000", x"000000", x"2004EB",
   x"820000", x"E0008A", x"3C04FE", x"820000", x"E000EA",
   x"3305B8", x"010000", x"B00022", x"490000", x"B00020",
   x"000000", x"000000", x"010001", x"B00021", x"000000",
   x"000000", x"010000", x"B00021", x"2005BA", x"490000",
   x"BA012C", x"010080", x"7000DF", x"3205C0", x"010002",
   x"C08127", x"8A0001", x"01FFFF", x"C0809B", x"890001",
   x"3305A5", x"400136", x"B0007B", x"01012C", x"B000A0",
   x"01001F", x"700137", x"0B0000", x"C000A0", x"870000",
   x"2004EB", x"1007E1", x"820000", x"E00088", x"3C04FE",
   x"4A0124", x"B80000", x"010080", x"7000DF", x"3205DA",
   x"010002", x"C080E2", x"8A0001", x"01FFFF", x"C0809B",
   x"880001", x"3305CF", x"000000", x"000000", x"2004EB",
   x"012000", x"7000DF", x"330684", x"010300", x"7000DF",
   x"E00099", x"3304F6", x"014000", x"7000DF", x"3205EF",
   x"490000", x"B00168", x"890001", x"2005F0", x"400168",
   x"0B0000", x"860000", x"018000", x"7000DF", x"33063C",
   x"820000", x"E0008A", x"3C04FE", x"820000", x"E00088",
   x"3805FE", x"4A016E", x"000000", x"20062E", x"820000",
   x"330603", x"40007C", x"000000", x"20062E", x"820000",
   x"E00081", x"330609", x"40016F", x"000000", x"20062E",
   x"820000", x"E00082", x"33060F", x"4A016E", x"000000",
   x"20062E", x"820000", x"E00083", x"330616", x"010001",
   x"B000C1", x"1007F3", x"20062E", x"820000", x"E00084",
   x"33061D", x"010002", x"B000C1", x"1007F3", x"20062E",
   x"820000", x"E00085", x"330624", x"010004", x"B000C1",
   x"1007F3", x"20062E", x"820000", x"E00086", x"33062B",
   x"010008", x"B000C1", x"1007F3", x"20062E", x"010010",
   x"B000C1", x"1007F3", x"B80000", x"010080", x"7000DF",
   x"320635", x"010002", x"C08168", x"8A0001", x"01FFFF",
   x"C0809B", x"880001", x"3305F5", x"000000", x"000000",
   x"2004EB", x"820000", x"E0008A", x"3C04FE", x"490000",
   x"BA016E", x"820000", x"E00088", x"3C0677", x"000000",
   x"820000", x"33064A", x"000000", x"000000", x"200677",
   x"820000", x"E00081", x"330652", x"40007C", x"B000C6",
   x"000000", x"10080B", x"200677", x"820000", x"E00082",
   x"330658", x"000000", x"000000", x"200677", x"820000",
   x"E00083", x"33065F", x"010001", x"B000C1", x"1007F3",
   x"200677", x"820000", x"E00084", x"330666", x"010002",
   x"B000C1", x"1007F3", x"200677", x"820000", x"E00085",
   x"33066D", x"010004", x"B000C1", x"1007F3", x"200677",
   x"820000", x"E00086", x"330674", x"010008", x"B000C1",
   x"1007F3", x"200677", x"010010", x"B000C1", x"1007F3",
   x"8A0001", x"010080", x"7000DF", x"32067D", x"010002",
   x"C08168", x"01FFFF", x"C0809B", x"890001", x"33063C",
   x"000000", x"000000", x"2004EB", x"1007E1", x"820000",
   x"E00088", x"3C04FE", x"4A0165", x"B80000", x"010080",
   x"7000DF", x"320690", x"010002", x"C080E2", x"8A0001",
   x"01FFFF", x"C0809B", x"880001", x"330685", x"000000",
   x"000000", x"2004EB", x"1007E1", x"820000", x"E00088",
   x"3C04FE", x"4A0154", x"B80000", x"010080", x"7000DF",
   x"3206A3", x"010002", x"C080E2", x"8A0001", x"01FFFF",
   x"C0809B", x"880001", x"330698", x"000000", x"000000",
   x"2004EB", x"012000", x"7000DF", x"3306F4", x"010300",
   x"7000DF", x"E00099", x"3304F6", x"014000", x"7000DF",
   x"3206B8", x"490000", x"B0015F", x"890001", x"2006B9",
   x"40015F", x"0B0000", x"860000", x"010002", x"70015F",
   x"3206C2", x"01C000", x"50015F", x"B000E0", x"2006C5",
   x"013000", x"50015F", x"B000E0", x"018000", x"7000DF",
   x"3306DE", x"010F00", x"7000E0", x"3304FE", x"000000",
   x"4000E0", x"100156", x"40009F", x"B80000", x"010080",
   x"7000DF", x"3206D7", x"010002", x"C0815F", x"010002",
   x"C080E0", x"01FFFF", x"C0809B", x"880001", x"3306C8",
   x"000000", x"000000", x"2004EB", x"010F00", x"7000E0",
   x"3304FE", x"490000", x"B0009E", x"4000E0", x"100143",
   x"010080", x"7000DF", x"3206ED", x"010002", x"C0815F",
   x"010002", x"C080E0", x"8A0001", x"01FFFF", x"C0809B",
   x"890001", x"3306DE", x"000000", x"000000", x"2004EB",
   x"1007E1", x"820000", x"E00088", x"3C04FE", x"4A015C",
   x"B80000", x"010080", x"7000DF", x"320700", x"010002",
   x"C080E2", x"8A0001", x"01FFFF", x"C0809B", x"880001",
   x"3306F5", x"000000", x"000000", x"2004EB", x"012000",
   x"7000DF", x"330755", x"010300", x"7000DF", x"E00099",
   x"3304F6", x"014000", x"7000DF", x"320715", x"490000",
   x"B0011F", x"890001", x"200716", x"40011F", x"0B0000",
   x"860000", x"B000D5", x"018000", x"7000DF", x"330738",
   x"01FFC0", x"7000D5", x"3304FE", x"000000", x"000000",
   x"100812", x"010003", x"E000D5", x"330728", x"4000D4",
   x"70008C", x"200729", x"4000D4", x"B80000", x"010080",
   x"7000DF", x"320731", x"010002", x"C0811F", x"010001",
   x"C080D5", x"01FFFF", x"C0809B", x"880001", x"33071C",
   x"000000", x"000000", x"2004EB", x"013602", x"E00139",
   x"320741", x"015A02", x"E00139", x"330506", x"01000F",
   x"E000D5", x"3C0506", x"01FFC0", x"7000D5", x"3304FE",
   x"490000", x"B000D3", x"10081B", x"010080", x"7000DF",
   x"32074E", x"010002", x"C0811F", x"010001", x"C080D5",
   x"01FFFF", x"C0809B", x"890001", x"330738", x"000000",
   x"000000", x"2004EB", x"1007E1", x"820000", x"E00088",
   x"3C04FE", x"4A011C", x"B80000", x"010080", x"7000DF",
   x"320761", x"010002", x"C080E2", x"8A0001", x"01FFFF",
   x"C0809B", x"880001", x"330756", x"000000", x"000000",
   x"2004EB", x"012000", x"7000DF", x"3307CE", x"014000",
   x"7000DF", x"320772", x"490000", x"B00103", x"890001",
   x"200773", x"400103", x"860000", x"012000", x"7000DF",
   x"3307CE", x"010300", x"7000DF", x"E0009A", x"3304F6",
   x"018000", x"7000DF", x"3307A4", x"800000", x"E000BA",
   x"3C04FE", x"400103", x"32078A", x"E00084", x"320790",
   x"E00084", x"320796", x"000000", x"000000", x"2004FE",
   x"100911", x"4000E4", x"B80000", x"4000E5", x"B80001",
   x"20079C", x"1008CA", x"010004", x"C080E4", x"010000",
   x"D080E5", x"200798", x"100911", x"1008E3", x"4000E6",
   x"B80000", x"4000E7", x"B80001", x"01FFFF", x"C0809B",
   x"000000", x"880002", x"33077E", x"000000", x"000000",
   x"2004EB", x"400103", x"3207AD", x"E00084", x"3207BB",
   x"E00088", x"3207B3", x"000000", x"000000", x"2004FE",
   x"100911", x"490000", x"B000E4", x"490001", x"B000E5",
   x"2007C7", x"100911", x"015A03", x"E00139", x"330506",
   x"000000", x"000000", x"100906", x"2007C7", x"015A03",
   x"E00139", x"330506", x"490000", x"B000E6", x"490001",
   x"B000E7", x"1008F0", x"010004", x"C080E4", x"010000",
   x"D080E5", x"01FFFF", x"C0809B", x"890002", x"3307A4",
   x"000000", x"000000", x"2004EB", x"1007E1", x"820000",
   x"E00088", x"3C04FE", x"4A0100", x"B80000", x"010080",
   x"7000DF", x"3207DA", x"010003", x"C080E2", x"8A0001",
   x"01FFFF", x"C0809B", x"880001", x"3307CF", x"000000",
   x"000000", x"2004EB", x"010300", x"7000DF", x"E00099",
   x"3304F6", x"018000", x"7000DF", x"330506", x"014000",
   x"7000DF", x"3207EF", x"490000", x"B000E2", x"890001",
   x"2007F0", x"4000E2", x"0B0000", x"860000", x"280000",
   x"010000", x"B000C5", x"40007C", x"B000C4", x"400070",
   x"7000C1", x"B000C3", x"400070", x"7000C1", x"B000C2",
   x"320800", x"4000C3", x"320809", x"4000C2", x"B000C3",
   x"40007C", x"E000C4", x"B000C5", x"E00170", x"3807FA",
   x"010020", x"50812C", x"4000C5", x"280000", x"40007C",
   x"E000C6", x"E0016F", x"38080B", x"000000", x"000000",
   x"280000", x"10088C", x"010006", x"10085C", x"4000D5",
   x"10086F", x"100897", x"B000D4", x"100893", x"280000",
   x"10088C", x"010004", x"10085C", x"01003F", x"10086F",
   x"100893", x"10088C", x"010005", x"10085C", x"4000D5",
   x"10086F", x"100848", x"10084E", x"4000D3", x"1008A8",
   x"100893", x"1008BB", x"10088C", x"010004", x"10085C",
   x"010000", x"10086F", x"100893", x"280000", x"010002",
   x"5080D2", x"280000", x"01FFFD", x"7080D2", x"280000",
   x"010001", x"5080D2", x"280000", x"01FFFE", x"7080D2",
   x"280000", x"330845", x"000000", x"000000", x"01FFFB",
   x"7080D2", x"280000", x"010004", x"5080D2", x"280000",
   x"010020", x"5080D2", x"280000", x"01FFDF", x"7080D2",
   x"280000", x"B0009E", x"01C022", x"100143", x"280000",
   x"01C022", x"100156", x"010008", x"70009F", x"280000",
   x"100833", x"10084E", x"100836", x"10084E", x"280000",
   x"B000A0", x"000000", x"000000", x"010004", x"7000A0",
   x"10083F", x"10084E", x"100857", x"010002", x"7000A0",
   x"10083F", x"10084E", x"100857", x"010001", x"7000A0",
   x"10083F", x"10084E", x"100857", x"280000", x"B000A0",
   x"010020", x"B000D6", x"000000", x"000000", x"4000A0",
   x"7000D6", x"10083F", x"10084E", x"4000D6", x"C00080",
   x"050000", x"B000D6", x"100833", x"10084E", x"100836",
   x"4000D6", x"330885", x"000000", x"000000", x"10084B",
   x"200886", x"100848", x"10084E", x"4000D6", x"330874",
   x"000000", x"000000", x"280000", x"010000", x"B000D2",
   x"10084E", x"010031", x"B000D2", x"10084E", x"280000",
   x"010000", x"B000D2", x"10084E", x"280000", x"B000A0",
   x"018000", x"B000D6", x"100857", x"100852", x"32089F",
   x"4000D6", x"5080A0", x"100857", x"4000D6", x"C00080",
   x"050000", x"B000D6", x"33089B", x"4000A0", x"000000",
   x"280000", x"B000A0", x"018000", x"B000D6", x"000000",
   x"000000", x"4000A0", x"7000D6", x"10083F", x"10084E",
   x"100857", x"4000D6", x"C00080", x"050000", x"B000D6",
   x"000000", x"3308AD", x"000000", x"000000", x"280000",
   x"01C350", x"B000A0", x"010011", x"B000D2", x"10084E",
   x"100852", x"3308C8", x"01FFFF", x"C080A0", x"3308C0",
   x"000000", x"000000", x"200506", x"100893", x"280000",
   x"01AA02", x"E000E8", x"3208D4", x"01AA02", x"B000E8",
   x"010000", x"B0007D", x"010003", x"10092F", x"100938",
   x"010000", x"10092F", x"B000E6", x"010000", x"10092F",
   x"060000", x"5080E6", x"010000", x"10092F", x"B000E7",
   x"010000", x"10092F", x"060000", x"5080E7", x"280000",
   x"010000", x"B0007D", x"0100AB", x"10092F", x"100938",
   x"010000", x"10092F", x"B000E6", x"010000", x"B000E7",
   x"01FFFF", x"B0007D", x"280000", x"01AA03", x"E000E8",
   x"3208FB", x"01AA03", x"B000E8", x"10094A", x"010000",
   x"B0007D", x"010002", x"10092F", x"100938", x"4000E6",
   x"10092F", x"4000E6", x"060000", x"10092F", x"4000E7",
   x"10092F", x"4000E7", x"060000", x"10092F", x"280000",
   x"10094A", x"010000", x"B0007D", x"0100D8", x"10092F",
   x"100938", x"010BB8", x"10091E", x"01AA01", x"B000E8",
   x"280000", x"01AA03", x"E000E8", x"320919", x"01FFFF",
   x"B0007D", x"01AA01", x"B000E8", x"280000", x"010005",
   x"10091E", x"01AA01", x"B000E8", x"280000", x"B0009C",
   x"01FFFF", x"B0007D", x"100940", x"700081", x"32092D",
   x"000000", x"010001", x"100450", x"01FFFF", x"C0809C",
   x"330921", x"000000", x"000000", x"200506", x"100951",
   x"280000", x"B0007E", x"000000", x"010002", x"70007D",
   x"330930", x"0100FF", x"70007E", x"B000E9", x"280000",
   x"4000E5", x"10092F", x"4000E4", x"060000", x"10092F",
   x"4000E4", x"10092F", x"280000", x"010000", x"B0007D",
   x"010005", x"10092F", x"010000", x"10092F", x"01FFFF",
   x"B0007D", x"4000E9", x"280000", x"010000", x"B0007D",
   x"010006", x"10092F", x"010001", x"B0007D", x"280000",
   x"010000", x"B0007D", x"010004", x"10092F", x"010001",
   x"B0007D", x"280000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"000000", x"000000", x"000000", x"000000", x"000000",
   x"00ABCD");

signal daddr: std_logic_vector(11 downto 0);

begin
   aetherhm2: process (clk)
   begin
      if (clk'event and clk = '1') then
         if (we = '1') then
            RAM(conv_integer(addr)) <= din;
         end if;
         daddr <= addr;
      end if; -- clk 
   end process;

   dout <= RAM(conv_integer(daddr));
end;
